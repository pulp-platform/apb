// Copyright (c) 2014 ETH Zurich, University of Bologna
//
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

// An APB4 (v2.0) interface
interface APB (
  parameter int unsigned AddrWidth = 32'd32,
  parameter int unsigned DataWidth = 32'd32,
  parameter int unsigned PselWidth = 32'd1
);
  localparam int unsigned StrbWidth = cf_math_pkg::ceil_div(DataWidth, 8);
  typedef logic [AddrWidth-1:0] addr_t;
  typedef logic [PselWidth-1:0] psel_t;
  typedef logic [DataWidth-1:0] data_t;
  typedef logic [StrbWidth-1:0] strb_t;

  addr_t          paddr;
  apb_pkg::prot_t pprot;
  psel_t          psel;
  logic           penable;
  logic           pwrite;
  data_t          pwdata;
  strb_t          pstrb;
  logic           pready;
  data_t          prdata;
  logic           pslverr;

  modport Master (
    output paddr, pprot, psel, penable, pwrite, pwdata, pstrb,
    input  pready, prdata, pslverr
  );

  modport Slave (
    input  paddr, pprot, psel, penable, pwrite, pwdata, pstrb,
    output pready, prdata, pslverr
  );

endinterface

// A clocked APB4 (v2.0) interface for use in design verification
interface APB_DV #(
  parameter int unsigned AddrWidth = 32'd32,
  parameter int unsigned DataWidth = 32'd32,
  parameter int unsigned PselWidth = 32'd1
) (
  input logic clk_i
);
  localparam int unsigned StrbWidth = cf_math_pkg::ceil_div(DataWidth, 8);
  typedef logic [AddrWidth-1:0] addr_t;
  typedef logic [PselWidth-1:0] psel_t;
  typedef logic [DataWidth-1:0] data_t;
  typedef logic [StrbWidth-1:0] strb_t;

  apb_pkg::addr_t paddr;
  apb_pkg::prot_t pprot;
  psel_t          psel;
  logic           penable;
  logic           pwrite;
  apb_pkg::data_t pwdata;
  apb_pkg::strb_t pstrb;
  logic           pready;
  apb_pkg::data_t prdata;
  logic           pslverr;

  modport Master (
    output paddr, pprot, psel, penable, pwrite, pwdata, pstrb,
    input  pready, prdata, pslverr
  );

  modport Slave (
    input  paddr, pprot, psel, penable, pwrite, pwdata, pstrb,
    output pready, prdata, pslverr
  );

endinterface
